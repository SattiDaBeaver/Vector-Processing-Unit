module mac_cell #(
    parameter DATA_WIDTH = 8,
    parameter ACC_WIDTH = 32
) (
    input  logic    in_a,
    input  logic    in_b
);
    
endmodule