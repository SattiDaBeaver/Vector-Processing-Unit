module tiny_fsm_control #(
    
) (

);

endmodule : tiny_fsm_control